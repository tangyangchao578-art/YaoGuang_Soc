//-----------------------------------------------------------------------------
// File: l3_cache_driver.sv
// Description: L3 Cache driver
// Author: YaoGuang SoC DV Team
// Date: 2026-01-18
//-----------------------------------------------------------------------------
`ifndef L3_CACHE_DRIVER_SV
`define L3_CACHE_DRIVER_SV

class l3_cache_driver extends uvm_driver#(l3_cache_transaction);
    `uvm_component_utils(l3_cache_driver)

    virtual l3_cache_if vif;
    l3_cache_config cfg;
    int transaction_count = 0;

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        if(!uvm_config_db#(virtual l3_cache_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("L3_CACHE_DRIVER", "Virtual interface not found")
        end
        cfg = l3_cache_config::type_id::create("cfg", this);
    endfunction

    task run_phase(uvm_phase phase);
        super.run_phase(phase);
        reset_driver();
        forever begin
            seq_item_port.get_next_item(req);
            drive_transaction(req);
            seq_item_port.item_done();
            transaction_count++;
        end
    endtask

    virtual task reset_driver();
        vif.valid <= 0;
        vif.ready <= 1;
        @(posedge vif.clk);
        #1;
    endtask

    virtual task drive_transaction(l3_cache_transaction tr);
        @(posedge vif.clk);
        vif.valid <= 1;
        vif.addr <= tr.addr;
        vif.data <= tr.data;
        vif.op <= tr.op;
        vif.id <= tr.id;
        vif.size <= tr.size;

        while(!vif.ready) begin
            @(posedge vif.clk);
            #0.1;
        end

        @(posedge vif.clk);
        vif.valid <= 0;
    endtask
endclass

`endif
