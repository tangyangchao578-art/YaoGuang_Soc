`ifndef DV_PKG_SVH
`define DV_PKG_SVH

package dv_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "dv_macros.svh"

`include "dv_config.svh"
`include "dv_sequence_item.svh"
`include "dv_sequence.svh"
`include "dv_driver.svh"
`include "dv_monitor.svh"
`include "dv_sequencer.svh"
`include "dv_agent.svh"
`include "dv_scoreboard.svh"
`include "dv_coverage.svh"
`include "dv_env.svh"

endpackage

`endif
